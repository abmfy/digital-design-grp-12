package util_func;
    function logic inside_range(int x, int a, int b);
        return a <= x && x < b;
    endfunction
endpackage